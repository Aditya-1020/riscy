/// instruciton cache
`timescale 1ps/1ps
`default_nettype none
`include "isa.v"

module icache (
    
);
    
endmodule